module i2c;







endmodule
